//////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX32_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: I0-I31 (32-bits each);  S (4-bit)
reg[31:0] I[31:0];
reg[4:0] S;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Y (32-bit)
wire[31:0] Y;
///////////////////////////////////////////////////////////////////////////////////

MUX32_32 myMUX(.I0(I[0]),.I1(I[1]),.I2(I[2]),.I3(I[3]),.I4(I[4]),.I5(I[5]),.I6(I[6]),.I7(I[7]),
.I8(I[8]),.I9(I[9]),.I_10(I[10]),.I_11(I[11]),.I_12(I[12]),.I_13(I[13]),.I_14(I[14]),.I_15(I[15]),
.I_16(I[16]),.I_17(I[17]),.I_18(I[18]),.I_19(I[19]),.I_20(I[20]),.I_21(I[21]),.I_22(I[22]),.I_23(I[23]),
.I_24(I[24]),.I_25(I[25]),.I_26(I[26]),.I_27(I[27]),.I_28(I[28]),.I_29(I[29]),.I_30(I[30]),.I_31(I[31]),.S(S),.Y(Y));

integer j;

initial begin

//////////////////////////////////////////////////////////////////////////////
// Initialize 32 input values
for (j = 0; j <= 31; j = j + 1) begin
  I[j] = (2**j)-1;
end
//////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////
//  Testing: All 5-bit S values 0 to 31
for (S=5'b00000; S <= 5'b11111; S = S + 5'b00001) begin
   $display("Testing: S=%b", S);
   #10;
   verifyEqual32(Y, I[S]);
   // You need this because the counter will reset to 0 otherwise
   if (S == 5'b11111) begin
    $display("All tests passed.");
    $stop;
   end
end
////////////////////////////////////////////////////////////////////////////////////////
  
end

endmodule